library verilog;
use verilog.vl_types.all;
entity CypherDetectorTB is
    port(
        d               : in     vl_logic
    );
end CypherDetectorTB;
