// qsys_files.v

// Generated using ACDS version 13.1 162 at 2023.01.02.08:22:51

`timescale 1 ps / 1 ps
module qsys_files (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
